module And_Gate_Data_Flow(a,b,y);
input a,b;
output y;
assign y = a&b;
endmodule
